`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:32:23 03/31/2015 
// Design Name: 
// Module Name:    piledArraySpliter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

/*
piledArr
{C3,B3,A3, C2,B2,A2, C1,B1,A1, C0,B0,A0}

piledArraySpliter

split into maximum four  arrays

*/
module piledArraySpliter
#(
parameter 



piledArrW=32
ArrL=32
)(
input 


    );


endmodule
